*TTL fanout calculation

.model Q1 npn Bf=50
Q11 2 1 0 Q1
Q12 1 5 4 Q1
R2 2 3 1.6K
R1 5 3 4K
Vcc 3 0 5
Vin 4 0 5

.subckt ttl out in c 0
Q21 out y 0 Q1
Q22 y z in Q1
R21 out c 1.6K
R11 z c 4K
.ends ttl

x1 out1 2 3 0 ttl
x2 out2 2 3 0 ttl
x3 out3 2 3 0 ttl
x4 out4 2 3 0 ttl
x5 out5 2 3 0 ttl
x6 out6 2 3 0 ttl
x7 out7 2 3 0 ttl
*x8 out8 2 3 0 ttl 		for 830 Vih

.dc Vin 0 5 0.05
.control
run
plot v(2) v(4)
.endc
.end