*TTL Inverter Transient Analysis

.model switch NPN (Bf=20)
Q1 2 1 4 switch
Q2 3 2 0 switch
R2 5 3 1.6k
R1 5 1 4k
Vcc 5 0 5
Vin 4 0 pulse(0 5 1ns 1ns 1ns 20us 40us)
c 3 0 1p
.tran 1ns 80us
.control
run
plot v(3) v(4)
.endc
.end
