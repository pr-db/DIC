*CMOS inverter

.model myPMOS PMOS (Vt0 = -1 Kp = 20u)
.model myNMOS NMOS (Vt0 = 0.8 Kp = 50u)

Vcc1 c1 0 5
Vcc2 c2 0 4
Vcc3 c3 0 3

Vin in 0 5


Mp1 out1 in c1 c1 myPMOS w=1.51u l=1u
Mn1 out1 in 0 0 myNMOS w=1u l=1u

Mp2 out2 in c2 c2 myPMOS w=1.51u l=1u
Mn2 out2 in 0 0 myNMOS w=1u l=1u

Mp3 out3 in c3 c3 myPMOS w=1.51u l=1u
Mn3 out3 in 0 0 myNMOS w=1u l=1u

.dc Vin 0 5 0.05
.control
run

plot V(in) V(out1) V(out2) V(out3)
.endc
.end
