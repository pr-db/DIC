*NMOS inverter

.model myNMOS NMOS(Vt0 =0.8 Kp = 20u)

Vin in 0 5
Vcc c 0 5

R1 c out1 100k
M1 out1 in 0 0 myNMOS w=2u l = 1u

R2 c out2 200k
M2 out2 in 0 0 myNMOS w=2u l = 1u

R3 c out3 300k
M3 out3 in 0 0 myNMOS w=2u l = 1u
.dc Vin 0 5 0.05
.control
run

Plot V(in) V(out1) V(out2) V(out3)
.endc
.end
