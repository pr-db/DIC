*RTL inverter fanout 

.model switch NPN Bf=20 

Q 2 1 0 switch
Rc 2 3 1k
Rb 4 1 10k
Vcc 3 0 5
Vin 4 0 5


.subckt rt1 out in c 0
q2 out y 0 switch
Rb1 in y 10k
Rc1 c out 1k
.ends Rt1 

X1 out1 2 3 0 Rt1
X2 out2 2 3 0 Rt1
X3 out3 2 3 0 Rt1
X4 out4 2 3 0 Rt1
X5 out5 2 3 0 Rt1
X6 out6 2 3 0 Rt1
X7 out7 2 3 0 Rt1
X8 out8 2 3 0 Rt1 

.dc Vin 0 5 0.05 

.control
run
plot V(2) V(4)
*plot V(out1)
.endc
.end
